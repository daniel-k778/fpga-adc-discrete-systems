// adc_subsystem.sv
//
// Wraps: XADC (VAUXP15/VAUXN15) + ready pulse + optional moving average + fixed-point mV scaler.
// Default scaling maps full-scale (FFFFh) ≈ 3300 (millivolts).
//
// Notes (per lab):
// - Channel: VAUXP15/VAUXN15 on Basys-3 JXADC (N2/N1). :contentReference[oaicite:6]{index=6}
// - XADC wizard: single-ended, continuous mode, ~1 MSPS, channel averaging enabled. :contentReference[oaicite:7]{index=7}
// - Extra moving-average improves effective resolution; reset causes "count-up" while window fills. :contentReference[oaicite:8]{index=8}
//
// Parameter guide:
//   AVG_POWER   = log2(window) for moving average (2^AVG_POWER samples). Set 0 to bypass averager.
//   AVG_WIDTH   = bit width carried through averager (typically 16).
//   SCALE_INT   / SCALE_SHIFT implement integer*value >> shift fixed-point scaling.
//
// Integrate: Instantiate here, wire vauxp15/vauxn15 from top pins/XDC, consume scaled/avg/raw.

module adc_subsystem #(
  parameter int unsigned AVG_POWER  = 12,   // 2^12 = 4096-sample moving average (set 0 to bypass)
  parameter int unsigned AVG_WIDTH  = 16,   // width of averaged output
  // Scale avg16 (0..65535) to millivolts (0..3300): scaled = (avg16 * 3300) >> 16
  parameter int unsigned SCALE_INT  = 3300,
  parameter int unsigned SCALE_SHIFT= 16
)(
  input  logic        clk,
  input  logic        reset,

  // XADC analog pins (Basys-3 JXADC: vauxp15=N2, vauxn15=N1) :contentReference[oaicite:9]{index=9}
  input  logic        vauxp15,
  input  logic        vauxn15,

  // Outputs
  output logic [15:0] raw16,       // raw 16b from XADC (top 12 bits hold conversion)
  output logic [15:0] raw12_hex,   // raw 12-bit value aligned to [15:4] for hex display
  output logic [15:0] avg16,       // averaged 16-bit (extra bits from averaging)
  output logic [15:0] scaled_mV,   // scaled to mV-like units (FFFFh ≈ 9999d)
  output logic        sample_pulse,// 1-cycle pulse when a new sample is captured
  output logic        busy,        // XADC busy
  output logic        eos          // end-of-sequence (single channel still toggles)
);

  // XADC wires
  localparam logic [6:0] CHANNEL_ADDR = 7'h1F; // XA4/AD15 (XADC4)
  logic        drdy, den;
  logic [15:0] do_out;

  // XADC instance (generated by Vivado IP wizard)
  xadc_wiz_0 XADC_INST (
    .di_in     (16'h0000),
    .daddr_in  (CHANNEL_ADDR),
    .den_in    (den),       // enable on EOC
    .dwe_in    (1'b0),
    .drdy_out  (drdy),      // data ready
    .do_out    (do_out),    // data
    .dclk_in   (clk),
    .reset_in  (reset),
    .vp_in     (1'b0),
    .vn_in     (1'b0),
    .vauxp15   (vauxp15),
    .vauxn15   (vauxn15),
    .channel_out(),         // unused
    .eoc_out   (den),       // use EOC to drive next read
    .alarm_out (),          // unused
    .eos_out   (eos),
    .busy_out  (busy)
  );

  // Edge-pulse on DRDY
  logic drdy_q;
  always_ff @(posedge clk) begin
    if (reset) drdy_q <= 1'b0;
    else       drdy_q <= drdy;
  end
  assign sample_pulse = (~drdy_q) & drdy;

  // Register the raw 16-bit word when DRDY fires
  always_ff @(posedge clk) begin
    if (reset) raw16 <= '0;
    else if (sample_pulse) raw16 <= do_out;
  end

  // Present the 12-bit result aligned to [15:4] for hex display compatibility
  assign raw12_hex = {raw16[15:4]};

  // Optional extra moving average (2^AVG_POWER); allow bypass if AVG_POWER==0
  // Din expects 16-bit; Q provides 16-bit averaged value.
  generate
    if (AVG_POWER == 0) begin : NO_AVG
      always_ff @(posedge clk) begin
        if (reset) avg16 <= '0;
        else if (sample_pulse) avg16 <= raw16;
      end
    end else begin : USE_AVG
      averager #(
        .power (AVG_POWER), // window length = 2^power
        .N     (AVG_WIDTH)  // width
      ) AVERAGER (
        .reset (reset),
        .clk   (clk),
        .EN    (sample_pulse),
        .Din   (raw16),
        .Q     (avg16)
      );
    end
  endgenerate

  // Fixed-point scaling to millivolts (FFFFh -> ~3300)
  always_ff @(posedge clk) begin
    if (reset) scaled_mV <= '0;
    else if (sample_pulse) scaled_mV <= (avg16 * SCALE_INT) >> SCALE_SHIFT;
  end

endmodule
